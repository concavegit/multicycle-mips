module cpu #(parameter instruction="mem/data.dat")(input clk);
endmodule
